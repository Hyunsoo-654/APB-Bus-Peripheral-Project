`timescale 1ns / 1ps

module FND_Periph(
    // global signals
    input  logic        PCLK,
    input  logic        PRESET,
    // APB Interface Signals
    input  logic [ 3:0] PADDR,
    input  logic        PWRITE,
    input  logic        PENABLE,
    input  logic [31:0] PWDATA,
    input  logic        PSEL,
    output logic [31:0] PRDATA,
    output logic        PREADY,
    output logic [ 3:0] fndCom,
    output logic [ 7:0] fndFont
);


    logic [13:0] number;

    APB_SlaveIntf_FND U_APB_SlaveInterf_FND (.*);


    fndController U_FNDCNTL(
        .clk(PCLK),
        .reset(PRESET),
        .number(number),
        .fnd_com(fndCom),
        .fnd_font(fndFont)
    );

endmodule


module APB_SlaveIntf_FND (
    // global signals
    input  logic        PCLK,
    input  logic        PRESET,
    // APB Interface Signals
    input  logic [ 3:0] PADDR,
    input  logic        PWRITE,
    input  logic        PENABLE,
    input  logic [31:0] PWDATA,
    input  logic        PSEL,
    output logic [31:0] PRDATA,
    output logic        PREADY,
    // Internal Port
    output logic [ 13:0] number
);

    logic [31:0] slv_reg0;

    assign number  = slv_reg0[13:0];

    always_ff @(posedge PCLK, posedge PRESET) begin
        if (PRESET) begin
            slv_reg0 <= 32'd0;
            PRDATA   <= 32'd0;
        end else begin
            PREADY <= 1'b0;
            if (PSEL && PENABLE) begin
                PREADY <= 1'b1;
                if (PWRITE) begin
                    case (PADDR[3:2])
                        2'd0: slv_reg0 <= PWDATA;
                    endcase
                end else begin
                    case (PADDR[3:2])
                        2'd0: PRDATA <= slv_reg0;
                    endcase
                end
            end
        end
    end
endmodule


module fndController (
    input  logic        clk,
    input  logic        reset,
    input  logic [13:0] number,
    output logic [ 3:0] fnd_com,
    output logic [ 7:0] fnd_font
);
    logic tick_1khz;
    logic [1:0] w_count;
    logic [3:0] w_digit;
    logic [3:0] w_digit_1;
    logic [3:0] w_digit_10;
    logic [3:0] w_digit_100;
    logic [3:0] w_digit_1000;

    clk_div_1khz U_clk_div_1khz (
        .clk(clk),
        .reset(reset),
        .tick_1khz(tick_1khz)
    );

    counter_2bit U_counter_2bit(
        .clk(clk),
        .reset(reset),
        .tick(tick_1khz),
        .count(w_count)
    );

    decoder_2x4 U_decoder_2x4 (
        .x(w_count),
        .y(fnd_com)
    );

    digitSplitter U_digitSplitter(
        .number(number),
        .digit_1(w_digit_1),
        .digit_10(w_digit_10),
        .digit_100(w_digit_100),
        .digit_1000(w_digit_1000)
    );

    mux_4x1 U_mux_4x1 (
        .digit_1(w_digit_1),
        .digit_10(w_digit_10),
        .digit_100(w_digit_100),
        .digit_1000(w_digit_1000),
        .sel(w_count),
        .bcd(w_digit)
    );

    BCDtoFND_Decoder U_BCDtoFND_Decoder(
        .bcd(w_digit),
        .fnd(fnd_font)
    );

endmodule


module clk_div_1khz (
    input  logic clk,
    input  logic reset,
    output logic tick_1khz
);

    logic [$clog2(100_000 - 1) : 0] div_counter;

    always_ff @(posedge clk, posedge reset) begin
        if (reset) begin
            div_counter <= 0;
            tick_1khz   <= 1'b0;
        end else begin
            if(div_counter == 100_000 - 1) begin // 100M -> 1hz, 1khz -> 100M - 1000
                div_counter <= 0;
                tick_1khz   <= 1'b1;
            end else begin
                div_counter <= div_counter + 1;
                tick_1khz   <= 1'b0;
            end
        end
    end

endmodule

module counter_2bit (
    input  logic       clk,
    input  logic       reset,
    input  logic       tick,
    output logic [1:0] count
);

    always_ff @(posedge clk, posedge reset) begin
        if (reset) begin
            count <= 0;
        end else begin
            if (tick) begin
                count <= count + 1;
            end
        end
    end

endmodule

module decoder_2x4 (
    input  logic [1:0] x,
    output logic [3:0] y
);
    always_comb begin 
        case (x)
            2'b00: y = 4'b1110 ;
            2'b01: y = 4'b1101 ;
            2'b10: y = 4'b1011 ;
            2'b11: y = 4'b0111 ;
            default: y = 4'b1111;
        endcase
    end
endmodule

module digitSplitter (
    input logic [13:0] number,
    output logic [3:0] digit_1,
    output logic [3:0] digit_10,
    output logic [3:0] digit_100,
    output logic [3:0] digit_1000
);

    assign digit_1 = number % 10;
    assign digit_10 = (number / 10) % 10;
    assign digit_100 = (number / 100) % 10;
    assign digit_1000 = (number / 1000) % 10;
    
endmodule

module mux_4x1 (
    input  logic [3:0] digit_1,
    input  logic [3:0] digit_10,
    input  logic [3:0] digit_100,
    input  logic [3:0] digit_1000,
    input  logic [1:0] sel,
    output logic [3:0] bcd
);

    always_comb begin
        case (sel)
            2'b00: bcd = digit_1;
            2'b01: bcd = digit_10;
            2'b10: bcd = digit_100;
            2'b11: bcd = digit_1000;
            default: bcd = 0;
        endcase
    end

endmodule

module BCDtoFND_Decoder (
    input  logic [3:0] bcd,
    output logic [7:0] fnd
);

    always_comb begin
        case (bcd)
            4'h0: fnd = 8'hc0;
            4'h1: fnd = 8'hf9;
            4'h2: fnd = 8'ha4;
            4'h3: fnd = 8'hb0;
            4'h4: fnd = 8'h99;
            4'h5: fnd = 8'h92;
            4'h6: fnd = 8'h82;
            4'h7: fnd = 8'hf8;
            4'h8: fnd = 8'h80;
            4'h9: fnd = 8'h90;
            4'ha: fnd = 8'h88;
            4'hb: fnd = 8'h83;
            4'hc: fnd = 8'hc6;
            4'hd: fnd = 8'ha1;
            4'he: fnd = 8'h86;
            4'hf: fnd = 8'h8e;
            default: fnd = 8'hff;
        endcase
    end

endmodule